//`include "mesi_isc_cpu_test.sv"

module mesi_isc_tb_wrp;
	mesi_isc_tb tb();
	cpu_sva_wrapper wrp();
endmodule
